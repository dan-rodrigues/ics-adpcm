`ifndef notes_vh
`define notes_vh

// 12 note scale encoded in 4bit values

`define NOTE_C  4'd0
`define NOTE_CS 4'd1
`define NOTE_D  4'd2
`define NOTE_DS 4'd3
`define NOTE_E  4'd4
`define NOTE_F  4'd5
`define NOTE_FS 4'd6
`define NOTE_G  4'd7
`define NOTE_GS 4'd8
`define NOTE_A  4'd9
`define NOTE_AS 4'd10
`define NOTE_B  4'd11

`define NOTE_UNDEFINED 4'd15

`endif
