`ifndef notes_vh
`define notes_vh

// 12 note scale encoded in 4bit values

`define NOTE_C  0
`define NOTE_CS 1
`define NOTE_D  2
`define NOTE_DS 3
`define NOTE_E  4
`define NOTE_F  5
`define NOTE_FS 6
`define NOTE_G  7
`define NOTE_GS 8
`define NOTE_A  9
`define NOTE_AS 10
`define NOTE_B  11

`define NOTE_UNDEFINED 15

`endif
